#include funciona por favor